`ifndef MEMORY_SVH
`define MEMORY_SVH

interface memory;
endinterface

`endif // MEMORY_SVH
