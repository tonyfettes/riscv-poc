`include "issue.svh"

module iq #(
  parameter SIZE = 3
) (
  input clock, reset,
  issue.iq issue,
);
endmodule
