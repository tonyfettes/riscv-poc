module core(
  input clock,
  input reset,
);
endmodule
