`include "defs.svh"

module ds #(
) (
);
endmodule
